module hazard(