library verilog;
use verilog.vl_types.all;
entity project1test is
end project1test;
