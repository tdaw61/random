library verilog;
use verilog.vl_types.all;
entity Project1_vlg_tst is
end Project1_vlg_tst;
