library verilog;
use verilog.vl_types.all;
entity fetchtest is
end fetchtest;
