library verilog;
use verilog.vl_types.all;
entity Test_regfile is
end Test_regfile;
