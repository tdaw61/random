library verilog;
use verilog.vl_types.all;
entity fetch_vlg_tst is
end fetch_vlg_tst;
