library verilog;
use verilog.vl_types.all;
entity proj2_vlg_tst is
end proj2_vlg_tst;
